module cpu;

endmodule
